--
--
--  This file is a part of JOP, the Java Optimized Processor
--
--  Copyright (C) 2001-2008, Martin Schoeberl (martin@jopdesign.com)
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--


--
--	bytecode.vhd
--
--	Show bytecode mnemonic in the simulation
--
--	Author: Martin Schoeberl	martin@jopdesign.com
--
--
--
--	2007-12-22	creation
--


library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bytecodectrl is

port (jinstr : in std_logic_vector(7 downto 0));
end bytecodectrl;

architecture sim of bytecodectrl is

	type bcval is (
			ctrl000,
ctrl001,
ctrl102,
ctrl103,
ctrl104,
ctrl105,
ctrl106,
ctrl107,
ctrl108,
ctrl109,
ctrl10A,
ctrl10B,
ctrl10C,
ctrl10D,
ctrl10E,
ctrl10F,
jopsys_clfz,
ctrl111,
ctrl112,
ctrl113,
ctrl114,
ctrl115,
ctrl116,
ctrl117,
ctrl118,
ctrl119,
ctrl11A,
ctrl11B,
ctrl11C,
ctrl11D,
ctrl11E,
ctrl11F,
ctrl120,
ctrl121,
ctrl122,
ctrl123,
ctrl124,
ctrl125,
ctrl126,
ctrl127,
ctrl128,
ctrl129,
ctrl12A,
ctrl12B,
ctrl12C,
ctrl12D,
ctrl12E,
jopsys_esl,
ctrl130,
ctrl131,
ctrl132,
ctrl133,
jopsys_noop,
ctrl135,
ctrl136,
ctrl137,
ctrl138,
ctrl139,
ctrl13A,
ctrl13B,
jopsys_cer,
ctrl13D,
jopsys_ceot,
jopsys_seot,
jopsys_ldrimm,
jopsys_cinit,
jopsys_strimm,
jopsys_subvimm, 
jopsys_subimm,
ctrl145,
ctrl146,
ctrl147,
jopsys_andimm,
ctrl149,
ctrl14A,
ctrl14B,
jopsys_orimm,
ctrl14D,
ctrl14E,
ctrl14F,
ctrl150,
ctrl151,
ctrl152,
ctrl153,
jopsys_sz,
ctrl155,
ctrl156,
ctrl157,
jopsys_jmpimm,
ctrl159,
ctrl15A,
ctrl15B,
jopsys_present,
ctrl15D,
ctrl15E,
ctrl15F,
ctrl160,
ctrl161,
ctrl162,
ctrl163,
ctrl164,
ctrl165,
ctrl166,
ctrl167,
ctrl168,
ctrl169,
ctrl16A,
ctrl16B,
ctrl16C,
ctrl16D,
ctrl16E,
ctrl16F,
ctrl170,
ctrl171,
ctrl172,
ctrl173,
ctrl174,
ctrl175,
ctrl176,
ctrl177,
jopsys_addimm,
ctrl179,
ctrl17A,
ctrl17B,
ctrl17C,
ctrl17D,
ctrl17E,
ctrl17F,
jopsys_ldrdir,
ctrl181,
jopsys_strdir,
ctrl183,
ctrl184,
ctrl185,
ctrl186,
ctrl187,
ctrl188,
ctrl189,
ctrl18A,
ctrl18B,
ctrl18C,
ctrl18D,
ctrl18E,
ctrl18F,
ctrl190,
ctrl191,
ctrl192,
ctrl193,
ctrl194,
ctrl195,
ctrl196,
ctrl197,
ctrl198,
ctrl199,
ctrl19A,
ctrl19B,
ctrl19C,
ctrl19D,
ctrl19E,
ctrl19F,
ctrl1A0,
ctrl1A1,
ctrl1A2,
ctrl1A3,
ctrl1A4,
ctrl1A5,
ctrl1A6,
ctrl1A7,
ctrl1A8,
ctrl1A9,
ctrl1AA,
ctrl1AB,
ctrl1AC,
ctrl1AD,
ctrl1AE,
ctrl1AF,
ctrl1B0,
ctrl1B1,
ctrl1B2,
ctrl1B3,
ctrl1B4,
ctrl1B5,
ctrl1B6,
ctrl1B7,
ctrl1B8,
ctrl1B9,
ctrl1BA,
ctrl1BB,
ctrl1BC,
ctrl1BD,
ctrl1BE,
ctrl1BF,
jopsys_ldind,
ctrl1C1,
jopsys_strind,
ctrl1C3,
ctrl1C4,
ctrl1C5,
ctrl1C6,
ctrl1C7,
jopsys_andind,
ctrl1C9,
ctrl1CA,
ctrl1CB,
jopsys_orind,
ctrl1CD,
ctrl1CE,
ctrl1CF,
ctrl1D0,
ctrl1D1,
ctrl1D2,
ctrl1D3,
ctrl1D4,
ctrl1D5,
ctrl1D6,
ctrl1D7,
jopsys_jmpind,
ctrl1D9,
ctrl1DA,
ctrl1DB,
ctrl1DC,
ctrl1DD,
ctrl1DE,
ctrl1DF,
jopsys_switchc,
ctrl1E1,
ctrl1E2,
ctrl1E3,
ctrl1E4,
ctrl1E5,
ctrl1E6,
ctrl1E7,
jopsys_datacall,
ctrl1E9,
ctrl1EA,
ctrl1EB,
jopsys_chkend,
ctrl1ED,
ctrl1EE,
ctrl1EF,
ctrl1F0,
ctrl1F1,
ctrl1F2,
ctrl1F3,
ctrl1F4,
ctrl1F5,
jopsys_ler,
jopsys_lsip,
jopsys_addind,
ctrl1F9,
jopsys_ssop,
jopsys_ssvop, 
ctrl1FC,
ctrl1FD,
ctrl1FE,
ctrl1FF
			--jopsys_ldrimm, jopsys_datacall
	);

	signal val : bcval;

begin

	val <= bcval'val(to_integer(unsigned(jinstr)));

end sim;
