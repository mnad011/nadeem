-- megafunction wizard: %RAM initializer%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTMEM_INIT 

-- ============================================================
-- File Name: xyz.vhd
-- Megafunction Name(s):
-- 			ALTMEM_INIT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Build 208 07/03/2011 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altmem_init CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" INIT_FILE="ctrl.mif" INIT_TO_ZERO="NO" NUMWORDS=16 PORT_ROM_DATA_READY="PORT_UNUSED" ROM_READ_LATENCY=1 WIDTH=1 WIDTHAD=4 clock dataout init init_busy ram_address ram_wren
--VERSION_BEGIN 11.0SP1 cbx_altmem_init 2011:07:03:21:05:55:SJ cbx_altsyncram 2011:07:03:21:05:55:SJ cbx_cycloneii 2011:07:03:21:05:55:SJ cbx_lpm_add_sub 2011:07:03:21:05:55:SJ cbx_lpm_compare 2011:07:03:21:05:55:SJ cbx_lpm_counter 2011:07:03:21:05:55:SJ cbx_lpm_decode 2011:07:03:21:05:55:SJ cbx_lpm_mux 2011:07:03:21:05:55:SJ cbx_mgl 2011:07:03:21:07:56:SJ cbx_stratix 2011:07:03:21:05:55:SJ cbx_stratixii 2011:07:03:21:05:55:SJ cbx_stratixiii 2011:07:03:21:05:55:SJ cbx_stratixv 2011:07:03:21:05:55:SJ cbx_util_mgl 2011:07:03:21:05:55:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsyncram 1 lpm_compare 2 lpm_counter 2 reg 8 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  xyz_meminit_bpl IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 init	:	IN  STD_LOGIC;
		 init_busy	:	OUT  STD_LOGIC;
		 ram_address	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 ram_wren	:	OUT  STD_LOGIC
	 ); 
 END xyz_meminit_bpl;

 ARCHITECTURE RTL OF xyz_meminit_bpl IS

	 SIGNAL  wire_int_rom_q_a	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 capture_init	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_addr	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_delay_addr_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_state_reg_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 state_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_state_reg_sclr	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 wire_state_reg_sload	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_lg_w_lg_w_q_range29w32w48w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_lg_w_q_range29w32w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_lg_w_q_range29w32w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_lg_w_q_range29w32w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_q_range3w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_q_range2w5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_q_range28w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_q_range29w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_lg_w_q_range40w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_q_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_q_range3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_q_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_q_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_reg_w_q_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_addr_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_addr_cmpr_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_wait_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_wait_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_gnd_vector	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_ctr_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_addr_ctr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_state_reg_w_lg_w_lg_w_q_range40w56w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wait_ctr_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wait_ctr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_rom_addr_state58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clken59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_init54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addrct_eq_numwords :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addrct_lt_numwords :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  clken	:	STD_LOGIC;
	 SIGNAL  dataout_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  done_state :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  idle_state :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  ram_write_state :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reset_state_machine :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rom_addr_state :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rom_data_capture_state :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  state_machine_clken :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  waitct_eq_latency :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  waitct_lt_latency :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTH_ECCSTATUS	:	NATURAL := 3;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone II";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(WIDTH_ECCSTATUS-1 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd_vector <= "0";
	wire_w_lg_clken59w(0) <= clken AND rom_data_capture_state(0);
	wire_w_lg_init54w(0) <= init OR capture_init(0);
	addrct_eq_numwords(0) <= wire_addr_cmpr_aeb;
	addrct_lt_numwords(0) <= wire_addr_cmpr_alb;
	clken <= '1';
	dataout <= dataout_w;
	dataout_w <= wire_int_rom_q_a;
	done_state(0) <= (wire_state_reg_w_lg_w_q_range3w13w(0) AND (NOT state_reg(0)));
	idle_state(0) <= (((NOT state_reg(2)) AND wire_state_reg_w_lg_w_q_range2w5w(0)) AND (NOT state_reg(0)));
	init_busy <= capture_init(0);
	ram_address <= delay_addr;
	ram_wren <= ram_write_state(0);
	ram_write_state(0) <= (((NOT state_reg(2)) AND state_reg(1)) AND state_reg(0));
	reset_state_machine(0) <= (ram_write_state(0) AND addrct_lt_numwords(0));
	rom_addr_state(0) <= (((NOT state_reg(2)) AND wire_state_reg_w_lg_w_q_range2w5w(0)) AND state_reg(0));
	rom_data_capture_state(0) <= (((NOT state_reg(2)) AND state_reg(1)) AND (NOT state_reg(0)));
	state_machine_clken(0) <= (clken AND ((idle_state(0) AND capture_init(0)) OR ((rom_data_capture_state(0) OR done_state(0)) OR (capture_init(0) AND (((NOT (rom_addr_state(0) AND waitct_lt_latency(0))) OR (rom_addr_state(0) AND waitct_eq_latency(0))) OR (ram_write_state(0) AND addrct_eq_numwords(0)))))));
	waitct_eq_latency(0) <= wire_wait_cmpr_aeb;
	waitct_lt_latency(0) <= wire_wait_cmpr_alb;
	int_rom :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "ctrl.mif",
		NUMWORDS_A => 16,
		OPERATION_MODE => "ROM",
		WIDTH_A => 1,
		WIDTHAD_A => 4,
		INTENDED_DEVICE_FAMILY => "Cyclone II"
	  )
	  PORT MAP ( 
		address_a => wire_addr_ctr_q,
		clock0 => clock,
		clocken0 => clken,
		q_a => wire_int_rom_q_a,
		rden_a => rom_data_capture_state(0)
	  );
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN capture_init(0) <= (wire_w_lg_init54w(0) AND (NOT done_state(0)));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_delay_addr_ena(0) = '1') THEN delay_addr(0) <= wire_addr_ctr_q(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_delay_addr_ena(1) = '1') THEN delay_addr(1) <= wire_addr_ctr_q(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_delay_addr_ena(2) = '1') THEN delay_addr(2) <= wire_addr_ctr_q(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_delay_addr_ena(3) = '1') THEN delay_addr(3) <= wire_addr_ctr_q(3);
			END IF;
		END IF;
	END PROCESS;
	loop0 : FOR i IN 0 TO 3 GENERATE
		wire_delay_addr_ena(i) <= wire_w_lg_clken59w(0);
	END GENERATE loop0;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (state_machine_clken(0) = '1') THEN 
				IF (wire_state_reg_sclr(0) = '1') THEN state_reg(0) <= '0';
				ELSIF (wire_state_reg_sload(0) = '1') THEN state_reg(0) <= '1';
				ELSE state_reg(0) <= wire_state_reg_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (state_machine_clken(0) = '1') THEN 
				IF (wire_state_reg_sclr(1) = '1') THEN state_reg(1) <= '0';
				ELSIF (wire_state_reg_sload(1) = '1') THEN state_reg(1) <= '1';
				ELSE state_reg(1) <= wire_state_reg_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (state_machine_clken(0) = '1') THEN 
				IF (wire_state_reg_sclr(2) = '1') THEN state_reg(2) <= '0';
				ELSIF (wire_state_reg_sload(2) = '1') THEN state_reg(2) <= '1';
				ELSE state_reg(2) <= wire_state_reg_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_state_reg_d <= ( wire_state_reg_w_lg_w_lg_w_lg_w_q_range29w32w48w49w & wire_state_reg_w_lg_w_lg_w_q_range29w32w43w & wire_state_reg_w_lg_w_lg_w_q_range29w32w33w);
	wire_state_reg_sclr <= ( reset_state_machine & reset_state_machine & "0");
	wire_state_reg_sload <= ( "0" & "0" & reset_state_machine);
	wire_state_reg_w_lg_w_lg_w_lg_w_q_range29w32w48w49w(0) <= wire_state_reg_w_lg_w_lg_w_q_range29w32w48w(0) AND wire_state_reg_w_q_range28w(0);
	wire_state_reg_w_lg_w_lg_w_q_range29w32w33w(0) <= wire_state_reg_w_lg_w_q_range29w32w(0) AND wire_state_reg_w_lg_w_q_range28w31w(0);
	wire_state_reg_w_lg_w_lg_w_q_range29w32w43w(0) <= wire_state_reg_w_lg_w_q_range29w32w(0) AND wire_state_reg_w_lg_w_q_range40w42w(0);
	wire_state_reg_w_lg_w_lg_w_q_range29w32w48w(0) <= wire_state_reg_w_lg_w_q_range29w32w(0) AND wire_state_reg_w_q_range40w(0);
	wire_state_reg_w_lg_w_q_range3w13w(0) <= wire_state_reg_w_q_range3w(0) AND wire_state_reg_w_lg_w_q_range2w5w(0);
	wire_state_reg_w_lg_w_q_range2w5w(0) <= NOT wire_state_reg_w_q_range2w(0);
	wire_state_reg_w_lg_w_q_range28w31w(0) <= NOT wire_state_reg_w_q_range28w(0);
	wire_state_reg_w_lg_w_q_range29w32w(0) <= NOT wire_state_reg_w_q_range29w(0);
	wire_state_reg_w_lg_w_q_range40w42w(0) <= wire_state_reg_w_q_range40w(0) XOR wire_state_reg_w_q_range28w(0);
	wire_state_reg_w_q_range2w(0) <= state_reg(1);
	wire_state_reg_w_q_range3w(0) <= state_reg(2);
	wire_state_reg_w_q_range28w(0) <= state_reg(0);
	wire_state_reg_w_q_range40w(0) <= state_reg(1);
	wire_state_reg_w_q_range29w(0) <= state_reg(2);
	wire_addr_cmpr_datab <= (OTHERS => '1');
	addr_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		aeb => wire_addr_cmpr_aeb,
		alb => wire_addr_cmpr_alb,
		dataa => delay_addr,
		datab => wire_addr_cmpr_datab
	  );
	wait_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 1
	  )
	  PORT MAP ( 
		aeb => wire_wait_cmpr_aeb,
		alb => wire_wait_cmpr_alb,
		dataa => wire_wait_ctr_q,
		datab => wire_gnd_vector
	  );
	wire_addr_ctr_sclr <= wire_state_reg_w_lg_w_lg_w_q_range40w56w57w(0);
	wire_state_reg_w_lg_w_lg_w_q_range40w56w57w(0) <= (NOT state_reg(1)) AND wire_state_reg_w_lg_w_q_range28w31w(0);
	addr_ctr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_modulus => 16,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 4
	  )
	  PORT MAP ( 
		clk_en => clken,
		clock => clock,
		cnt_en => ram_write_state(0),
		q => wire_addr_ctr_q,
		sclr => wire_addr_ctr_sclr
	  );
	wire_wait_ctr_sclr <= wire_w_lg_rom_addr_state58w(0);
	wire_w_lg_rom_addr_state58w(0) <= NOT rom_addr_state(0);
	wait_ctr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_modulus => 1,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 1
	  )
	  PORT MAP ( 
		clk_en => clken,
		clock => clock,
		cnt_en => rom_addr_state(0),
		q => wire_wait_ctr_q,
		sclr => wire_wait_ctr_sclr
	  );

 END RTL; --xyz_meminit_bpl
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY xyz IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		init		: IN STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		init_busy		: OUT STD_LOGIC ;
		ram_address		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		ram_wren		: OUT STD_LOGIC 
	);
END xyz;


ARCHITECTURE RTL OF xyz IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC ;



	COMPONENT xyz_meminit_bpl
	PORT (
			clock	: IN STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			init	: IN STD_LOGIC ;
			init_busy	: OUT STD_LOGIC ;
			ram_address	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			ram_wren	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(0 DOWNTO 0);
	init_busy    <= sub_wire1;
	ram_address    <= sub_wire2(3 DOWNTO 0);
	ram_wren    <= sub_wire3;

	xyz_meminit_bpl_component : xyz_meminit_bpl
	PORT MAP (
		clock => clock,
		init => init,
		dataout => sub_wire0,
		init_busy => sub_wire1,
		ram_address => sub_wire2,
		ram_wren => sub_wire3
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: INIT_FILE STRING "ctrl.mif"
-- Retrieval info: CONSTANT: INIT_TO_ZERO STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmem_init"
-- Retrieval info: CONSTANT: NUMWORDS NUMERIC "16"
-- Retrieval info: CONSTANT: PORT_ROM_DATA_READY STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: ROM_READ_LATENCY NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTHAD NUMERIC "4"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataout 0 0 1 0 OUTPUT NODEFVAL "dataout[0..0]"
-- Retrieval info: CONNECT: dataout 0 0 1 0 @dataout 0 0 1 0
-- Retrieval info: USED_PORT: init 0 0 0 0 INPUT NODEFVAL "init"
-- Retrieval info: CONNECT: @init 0 0 0 0 init 0 0 0 0
-- Retrieval info: USED_PORT: init_busy 0 0 0 0 OUTPUT NODEFVAL "init_busy"
-- Retrieval info: CONNECT: init_busy 0 0 0 0 @init_busy 0 0 0 0
-- Retrieval info: USED_PORT: ram_address 0 0 4 0 OUTPUT NODEFVAL "ram_address[3..0]"
-- Retrieval info: CONNECT: ram_address 0 0 4 0 @ram_address 0 0 4 0
-- Retrieval info: USED_PORT: ram_wren 0 0 0 0 OUTPUT NODEFVAL "ram_wren"
-- Retrieval info: CONNECT: ram_wren 0 0 0 0 @ram_wren 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL xyz.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
